module axi2ahb #(
    // Width of ID for for write address, write data, read address and read data
    parameter integer AXI_ID_WIDTH   = 1,
    // Width of S_AXI data bus
    parameter integer AXI_DATA_WIDTH = 32,
    // Width of S_AXI address bus
    parameter integer AXI_ADDR_WIDTH = 8
) (
    // Global Clock Signal
    input  wire                            ACLK,
    // Global Reset Signal. This Signal                        is Active LOW
    input  wire                            ARESETN,
    // ==========================================================
    // Write address                                                       channel
    // ==========================================================
    // Write Address ID
    input  wire [      AXI_ID_WIDTH-1 : 0] AWID,
    // Write address
    input  wire [    AXI_ADDR_WIDTH-1 : 0] AWADDR,
    // Burst length. The burst length gives the exact number of transfers in a burst
    input  wire [                   7 : 0] AWLEN,
    // Burst size. This signal indicates the size of each transfer in the burst
    input  wire [                   2 : 0] AWSIZE,
    // Burst type. The burst type and the size information,
    // determine how the address for each transfer within the burst is calculated.
    input  wire [                   1 : 0] AWBURST,
    // Write address valid. This signal indicates that
    // the channel is signaling valid write address and
    // control information.
    input  wire                            AWVALID,
    // Write address ready. This signal indicates that
    // the slave is ready to accept an address and associated
    // control signals.
    output wire                            AWREADY,
    // ==========================================================
    // Write data channel
    // ==========================================================
    // Write Data
    input  wire [    AXI_DATA_WIDTH-1 : 0] WDATA,
    // Write strobes. This signal indicates which byte
    // lanes hold valid data. There is one write strobe
    // bit for each eight bits of the write data bus.
    input  wire [(AXI_DATA_WIDTH/8)-1 : 0] WSTRB,
    // Write last. This signal indicates the last transfer
    // in a write burst.
    input  wire                            WLAST,
    // Write valid. This signal indicates that valid write
    // data and strobes are available.
    input  wire                            WVALID,
    // Write ready. This signal indicates that the slave
    // can accept the write data.
    output wire                            WREADY,
    // ==========================================================
    // Write response channel
    // ==========================================================
    // Response ID tag. This signal is the ID tag of the
    // write response.
    output wire [      AXI_ID_WIDTH-1 : 0] BID,
    // Write response. This signal indicates the status
    // of the write transaction.
    output wire [                   1 : 0] BRESP,
    // Write response valid. This signal indicates that the
    // channel is signaling a valid write response.
    output wire                            BVALID,
    // Response ready. This signal indicates that the master
    // can accept a write response.
    input  wire                            BREADY,
    // ==========================================================
    // Read address channel
    // ==========================================================
    // Read address ID. This signal is the identification
    // tag for the read address group of signals.
    input  wire [      AXI_ID_WIDTH-1 : 0] ARID,
    // Read address. This signal indicates the initial
    // address of a read burst transaction.
    input  wire [    AXI_ADDR_WIDTH-1 : 0] ARADDR,
    // Burst length. The burst length gives the exact number of transfers in a burst
    input  wire [                   7 : 0] ARLEN,
    // Burst size. This signal indicates the size of each transfer in the burst
    input  wire [                   2 : 0] ARSIZE,
    // Burst type. The burst type and the size information,
    // determine how the address for each transfer within the burst is calculated.
    input  wire [                   1 : 0] ARBURST,
    // Write address valid. This signal indicates that
    // the channel is signaling valid read address and
    // control information.
    input  wire                            ARVALID,
    // Read address ready. This signal indicates that
    // the slave is ready to accept an address and associated
    // control signals.
    output wire                            ARREADY,
    // ==========================================================
    // Read data channel
    // ==========================================================
    // Read ID tag. This signal is the identification tag
    // for the read data group of signals generated by the slave.
    output wire [      AXI_ID_WIDTH-1 : 0] RID,
    // Read Data
    output wire [    AXI_DATA_WIDTH-1 : 0] RDATA,
    // Read response. This signal indicates the status of
    // the read transfer.
    output wire [                   1 : 0] RRESP,
    // Read last. This signal indicates the last transfer
    // in a read burst.
    output wire                            RLAST,
    // Read valid. This signal indicates that the channel
    // is signaling the required read data.
    output wire                            RVALID,
    // Read ready. This signal indicates that the master can
    // accept the read data and response information.
    input  wire                            RREADY,
    // ==========================================================
    // AHB Master Interface
    // ==========================================================
    output wire [      AXI_ADDR_WIDTH-1:0] HADDR,
    output wire [                     2:0] HBURST,
    output wire [                     2:0] HSIZE,
    output wire [                     1:0] HTRANS,
    output wire                            HWRITE,
    output wire [      AXI_DATA_WIDTH-1:0] HWDATA,
    input  wire                            HREADY,
    input  wire [      AXI_DATA_WIDTH-1:0] HRDATA
);

    wire [    AXI_ID_WIDTH-1:0] cmd_id;
    wire                        cmd_read;
    wire                        cmd_write;
    wire [AXI_ADDR_WIDTH-1 : 0] cmd_start_addr;
    wire [                 7:0] cmd_transfer_len;
    wire [                 1:0] cmd_burst_type;
    wire                        cmd_error;
    wire                        ctrl_cmd_valid;
    wire                        ctrl_cmd_ready;

    wire                        ctrl_read_ready;
    wire                        ctrl_read_valid;
    wire                        ctrl_read_last;

    wire                        ctrl_write_ready;
    wire                        ctrl_write_valid;
    wire                        ctrl_write_last;

    axi2ahb_cmd #(
        .AXI_ID_WIDTH  (AXI_ID_WIDTH),
        .AXI_ADDR_WIDTH(AXI_ADDR_WIDTH)
    ) bridge_cmd (
        .ACLK              (ACLK),
        .ARESETN           (ARESETN),
        // AXI Write address channel
        .AWID              (AWID),
        .AWADDR            (AWADDR),
        .AWLEN             (AWLEN),
        .AWSIZE            (AWSIZE),
        .AWBURST           (AWBURST),
        .AWVALID           (AWVALID),
        .AWREADY           (AWREADY),
        // AXI Read address channel
        .ARID              (ARID),
        .ARADDR            (ARADDR),
        .ARLEN             (ARLEN),
        .ARSIZE            (ARSIZE),
        .ARBURST           (ARBURST),
        .ARVALID           (ARVALID),
        .ARREADY           (ARREADY),
        // CMD dispatch interface
        .cmd_id_o          (cmd_id),
        .cmd_read_o        (cmd_read),
        .cmd_write_o       (cmd_write),
        .cmd_start_addr_o  (cmd_start_addr),
        .cmd_transfer_len_o(cmd_transfer_len),
        .cmd_burst_type_o  (cmd_burst_type),
        .cmd_error_o       (cmd_error),
        .ctrl_cmd_valid_o  (ctrl_cmd_valid),
        .ctrl_cmd_ready_i  (ctrl_cmd_ready)
    );

    axi2ahb_ctrl #(
        .AXI_ADDR_WIDTH(AXI_ADDR_WIDTH)
    ) bridge_ctrl (
        .ACLK              (ACLK),
        .ARESETN           (ARESETN),
        .HADDR             (HADDR),
        .HBURST            (HBURST),
        .HSIZE             (HSIZE),
        .HTRANS            (HTRANS),
        .HREADY            (HREADY),
        .HWRITE            (HWRITE),
        // CMD dispatch interface
        .cmd_read_i        (cmd_read),
        .cmd_write_i       (cmd_write),
        .cmd_start_addr_i  (cmd_start_addr),
        .cmd_transfer_len_i(cmd_transfer_len),
        .cmd_burst_type_i  (cmd_burst_type),
        .ctrl_cmd_valid_i  (ctrl_cmd_valid),
        .ctrl_cmd_ready_o  (ctrl_cmd_ready),
        // Ready-Write control interface
        .ctrl_rdata_ready_i(ctrl_rdata_ready),
        .ctrl_rdata_valid_o(ctrl_rdata_valid),
        .ctrl_rdata_last_o (ctrl_rdata_last),
        .ctrl_wdata_last_i (ctrl_wdata_last),
        .ctrl_wdata_ready_i(ctrl_wdata_ready),
        .ctrl_wdata_valid_o(ctrl_wdata_valid)
    );


    axi2ahb_wdata #(
        .AXI_ID_WIDTH  (AXI_ID_WIDTH),
        .AXI_DATA_WIDTH(AXI_DATA_WIDTH)
    ) bridge_wdata (
        .ACLK(ACLK),
        .ARESETN(ARESETN),
        .WDATA(WDATA),
        .WSTRB(WSTRB),
        .WLAST(WLAST),
        .WVALID(WVALID),
        .WREADY(WREADY),
        .BID(BID),
        .BRESP(BRESP),
        .BVALID(BVALID),
        .BREADY(BREADY),
        .HWDATA(HWDATA),
        .HREADY(HREADY),
        .cmd_id_i(cmd_id),
        .ctrl_wdata_last_o(ctrl_wdata_last),
        .ctrl_wdata_valid_i(ctrl_wdata_valid),
        .ctrl_wdata_ready_o(ctrl_wdata_ready)
    );


endmodule
